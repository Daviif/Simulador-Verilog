module alu_control(
    input logic [1:0] aluOp,
    input logic [2:0] funct3,
    input logic funct7,
    output logic [2:0] alu_control
);
    

endmodule
module imm_gen(
    input logic [31:0] instrucao,
    output logic [31:0] immediate
);

endmodule